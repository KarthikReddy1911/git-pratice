package pkg;
`include "transaction.sv"
`include "generator.sv"
`include "driver.sv"
`include "monitor.sv"
`include "refernce_model.sv"
`include "scoreboard.sv"
`include "environment.sv"
`include "test.sv"
endpackage
